module my_buffer (A, B);
  input A;
  output B;
  assign B=A;
endmodule
